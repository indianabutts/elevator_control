/// Button Panel Module for Hallway Control
// Has Up and Down and Illuminates the Direction when
// Ack is received from the Building Controller
// Will also Exclude the unneccessary button in the
// case of top and bottom floor

module button_hall(
);