

module top()

  buidling_dispatcher DISPATCH(.*);
   a
   


endmodule // top
