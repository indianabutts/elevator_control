//Global Parameters File
//To make it easy to change variables across the design

module global_parameters();

`define FLOOR_COUNT 7


endmodule; // global_parameters
