/// Building Controller
/// Handles the inputs from the Hallway buttons
/// and determines the best of the two elevators to
/// dispatch the request to
`timescale 1ns/1ps
module building_controller (
			    );
   

endmodule
